module estados ( 
	reset,
	x1,
	clk,
	z
	) ;

input  reset;
input [1:0] x1;
input  clk;
inout  z;
